
interface DecodedInsttruction ();

	wire test;

endinterface
